entity sim is end entity sim;

architecture sim of sim is
    component challenge0_sim is end component;

begin
    challenge0_sim_inst: challenge0_sim;
end architecture sim;

