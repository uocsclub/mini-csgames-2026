entity sim is end entity sim;

architecture sim of sim is
    component challenge0_sim is end component;
    component challenge1_sim is end component;
    component challenge2_sim is end component;

begin
    -- challenge0_sim_inst: challenge0_sim;
    -- challenge1_sim_inst: challenge1_sim;
    challenge2_sim_inst: challenge2_sim;
end architecture sim;

